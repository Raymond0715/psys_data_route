`define SIM
