//`define SIM_BD
