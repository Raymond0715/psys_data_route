`define SIM_BD
