`define DROUTE_SIM
